module main

#flag wasm32_emscripten --embed-file @DIR/resources/Graduate-Regular.ttf@/resources/Graduate-Regular.ttf
#flag wasm32_emscripten --embed-file @DIR/resources/player.png@/resources/player.png
#flag wasm32_emscripten --embed-file @DIR/resources/enemy.png@/resources/enemy.png
#flag wasm32_emscripten --embed-file @DIR/resources/water.png@/resources/water.png
#flag wasm32_emscripten --embed-file @DIR/resources/land.png@/resources/land.png
#flag wasm32_emscripten --embed-file @DIR/resources/ball.png@/resources/ball.png
